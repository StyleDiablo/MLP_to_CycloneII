library verilog;
use verilog.vl_types.all;
entity cyNet_vlg_vec_tst is
end cyNet_vlg_vec_tst;
