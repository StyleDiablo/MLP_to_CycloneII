library verilog;
use verilog.vl_types.all;
entity top_sim is
end top_sim;
